module riscv_pc ();
endmodule