library verilog;
use verilog.vl_types.all;
entity riscv_datapath is
    generic(
        width           : integer := 64;
        MXLEN           : integer := 64
    );
    port(
        i_riscv_datapath_clk: in     vl_logic;
        i_riscv_datapath_rst: in     vl_logic;
        i_riscv_datapath_stallpc: in     vl_logic;
        o_riscv_datapath_pc: out    vl_logic_vector;
        i_riscv_datapath_inst: in     vl_logic_vector(31 downto 0);
        i_riscv_datapath_flush_fd: in     vl_logic;
        i_riscv_datapath_stall_fd: in     vl_logic;
        i_riscv_datapath_immsrc: in     vl_logic_vector(2 downto 0);
        o_riscv_datapath_opcode: out    vl_logic_vector(6 downto 0);
        o_riscv_datapath_func3: out    vl_logic_vector(2 downto 0);
        o_riscv_datapath_func7_5: out    vl_logic;
        o_riscv_datapath_func7_0: out    vl_logic;
        o_riscv_datapath_rs1addr_d: out    vl_logic_vector(4 downto 0);
        o_riscv_datapath_rs2addr_d: out    vl_logic_vector(4 downto 0);
        i_riscv_datapath_regw: in     vl_logic;
        i_riscv_datapath_jump: in     vl_logic;
        i_riscv_datapath_asel: in     vl_logic;
        i_riscv_datapath_bsel: in     vl_logic;
        i_riscv_datapath_memw: in     vl_logic;
        i_riscv_datapath_memr: in     vl_logic;
        i_riscv_datapath_storesrc: in     vl_logic_vector(1 downto 0);
        i_riscv_datapath_resultsrc: in     vl_logic_vector(1 downto 0);
        i_riscv_datapath_bcond: in     vl_logic_vector(3 downto 0);
        i_riscv_datapath_memext: in     vl_logic_vector(2 downto 0);
        i_riscv_datapath_aluctrl: in     vl_logic_vector(5 downto 0);
        i_riscv_datapath_mulctrl: in     vl_logic_vector(3 downto 0);
        i_riscv_datapath_divctrl: in     vl_logic_vector(3 downto 0);
        i_riscv_datapath_funcsel: in     vl_logic_vector(1 downto 0);
        i_riscv_datapath_flush_de: in     vl_logic;
        i_riscv_datapath_fwda: in     vl_logic_vector(1 downto 0);
        i_riscv_datapath_fwdb: in     vl_logic_vector(1 downto 0);
        o_riscv_datapath_icu_valid_e: out    vl_logic;
        o_riscv_datapath_pcsrc_e: out    vl_logic;
        o_riscv_datapath_rs1addr_e: out    vl_logic_vector(4 downto 0);
        o_riscv_datapath_rs2addr_e: out    vl_logic_vector(4 downto 0);
        o_riscv_datapath_rdaddr_e: out    vl_logic_vector(4 downto 0);
        o_riscv_datapath_resultsrc_e: out    vl_logic_vector(1 downto 0);
        o_riscv_datapath_opcode_m: out    vl_logic_vector(6 downto 0);
        o_datapath_div_en: out    vl_logic;
        o_datapath_mul_en: out    vl_logic;
        i_riscv_datapath_dm_rdata: in     vl_logic_vector;
        o_riscv_datapath_rdaddr_m: out    vl_logic_vector(4 downto 0);
        o_riscv_datapath_memw_e: out    vl_logic;
        o_riscv_datapath_memr_e: out    vl_logic;
        o_riscv_datapath_storesrc_m: out    vl_logic_vector(1 downto 0);
        o_riscv_datapath_memodata_addr: out    vl_logic_vector;
        o_riscv_datapath_storedata_m: out    vl_logic_vector;
        o_riscv_datapath_regw_m: out    vl_logic;
        o_riscv_datapath_regw_wb: out    vl_logic;
        o_riscv_datapath_rdaddr_wb: out    vl_logic_vector(4 downto 0);
        i_riscv_datapath_stall_de: in     vl_logic;
        i_riscv_datapath_stall_em: in     vl_logic;
        i_riscv_datapath_stall_mw: in     vl_logic;
        i_riscv_datapath_illgalinst_cu_de: in     vl_logic;
        i_riscv_datapath_csrop_cu_de: in     vl_logic_vector(2 downto 0);
        i_riscv_datapath_iscsr_cu_de: in     vl_logic;
        i_riscv_datapath_ecallu_cu_de: in     vl_logic;
        i_riscv_datapath_ecalls_cu_de: in     vl_logic;
        i_riscv_datapath_ecallm_cu_de: in     vl_logic;
        i_riscv_datapath_immreg_cu_de: in     vl_logic;
        o_riscv_datapath_rs1_fd_cu: out    vl_logic_vector(4 downto 0);
        o_riscv_datapath_constimm12_fd_cu: out    vl_logic_vector(11 downto 0);
        i_riscv_core_timerinterupt: in     vl_logic;
        i_riscv_core_externalinterupt: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width : constant is 1;
    attribute mti_svvh_generic_type of MXLEN : constant is 1;
end riscv_datapath;
