module riscv_divider (
input  logic signed [63:0]   i_riscv_div_rs1data,
input  logic signed [63:0]   i_riscv_div_rs2data,
input  logic        [2:0]    i_riscv_div_divctrl,
output logic signed [63:0]   o_riscv_div_product
);



endmodule
