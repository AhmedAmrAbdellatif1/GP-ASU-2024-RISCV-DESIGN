//salam allikom 
//bgrab bas
