library verilog;
use verilog.vl_types.all;
entity riscv_de_ppreg is
    generic(
        width           : integer := 64
    );
    port(
        i_riscv_de_clk  : in     vl_logic;
        i_riscv_de_rst  : in     vl_logic;
        i_riscv_de_flush: in     vl_logic;
        i_riscv_de_en   : in     vl_logic;
        i_riscv_de_pc_d : in     vl_logic_vector(63 downto 0);
        i_riscv_de_rs1addr_d: in     vl_logic_vector(4 downto 0);
        i_riscv_de_rs1data_d: in     vl_logic_vector(63 downto 0);
        i_riscv_de_rs2data_d: in     vl_logic_vector(63 downto 0);
        i_riscv_de_rs2addr_d: in     vl_logic_vector(4 downto 0);
        i_riscv_de_rdaddr_d: in     vl_logic_vector(4 downto 0);
        i_riscv_de_extendedimm_d: in     vl_logic_vector(63 downto 0);
        i_riscv_de_b_condition_d: in     vl_logic_vector(3 downto 0);
        i_riscv_de_oprnd2sel_d: in     vl_logic;
        i_riscv_de_storesrc_d: in     vl_logic_vector(1 downto 0);
        i_riscv_de_alucontrol_d: in     vl_logic_vector(5 downto 0);
        i_riscv_de_mulctrl_d: in     vl_logic_vector(3 downto 0);
        i_riscv_de_divctrl_d: in     vl_logic_vector(3 downto 0);
        i_riscv_de_funcsel_d: in     vl_logic_vector(1 downto 0);
        i_riscv_de_oprnd1sel_d: in     vl_logic;
        i_riscv_de_memwrite_d: in     vl_logic;
        i_riscv_de_memread_d: in     vl_logic;
        i_riscv_de_memext_d: in     vl_logic_vector(2 downto 0);
        i_riscv_de_resultsrc_d: in     vl_logic_vector(1 downto 0);
        i_riscv_de_regwrite_d: in     vl_logic;
        i_riscv_de_jump_d: in     vl_logic;
        i_riscv_de_pcplus4_d: in     vl_logic_vector(63 downto 0);
        i_riscv_de_opcode_d: in     vl_logic_vector(6 downto 0);
        o_riscv_de_pc_e : out    vl_logic_vector(63 downto 0);
        o_riscv_de_pcplus4_e: out    vl_logic_vector(63 downto 0);
        o_riscv_de_rs1addr_e: out    vl_logic_vector(4 downto 0);
        o_riscv_de_rs1data_e: out    vl_logic_vector(63 downto 0);
        o_riscv_de_rs2data_e: out    vl_logic_vector(63 downto 0);
        o_riscv_de_rs2addr_e: out    vl_logic_vector(4 downto 0);
        o_riscv_de_rdaddr_e: out    vl_logic_vector(4 downto 0);
        o_riscv_de_extendedimm_e: out    vl_logic_vector(63 downto 0);
        o_riscv_de_b_condition_e: out    vl_logic_vector(3 downto 0);
        o_riscv_de_oprnd2sel_e: out    vl_logic;
        o_riscv_de_storesrc_e: out    vl_logic_vector(1 downto 0);
        o_riscv_de_alucontrol_e: out    vl_logic_vector(5 downto 0);
        o_riscv_de_mulctrl_e: out    vl_logic_vector(3 downto 0);
        o_riscv_de_divctrl_e: out    vl_logic_vector(3 downto 0);
        o_riscv_de_funcsel_e: out    vl_logic_vector(1 downto 0);
        o_riscv_de_oprnd1sel_e: out    vl_logic;
        o_riscv_de_memwrite_e: out    vl_logic;
        o_riscv_de_memread_e: out    vl_logic;
        o_riscv_de_memext_e: out    vl_logic_vector(2 downto 0);
        o_riscv_de_resultsrc_e: out    vl_logic_vector(1 downto 0);
        o_riscv_de_regwrite_e: out    vl_logic;
        o_riscv_de_jump_e: out    vl_logic;
        o_riscv_de_opcode_e: out    vl_logic_vector(6 downto 0);
        i_riscv_de_ecall_m_d: in     vl_logic;
        i_riscv_de_csraddress_d: in     vl_logic_vector(11 downto 0);
        i_riscv_de_illegal_inst_d: in     vl_logic;
        i_riscv_de_iscsr_d: in     vl_logic;
        i_riscv_de_csrop_d: in     vl_logic_vector(2 downto 0);
        i_riscv_de_immreg_d: in     vl_logic;
        i_riscv_de_immzeroextend_d: in     vl_logic_vector;
        o_riscv_de_ecall_m_e: out    vl_logic;
        o_riscv_de_csraddress_e: out    vl_logic_vector(11 downto 0);
        o_riscv_de_illegal_inst_e: out    vl_logic;
        o_riscv_de_iscsr_e: out    vl_logic;
        o_riscv_de_csrop_e: out    vl_logic_vector(2 downto 0);
        o_riscv_de_immreg_e: out    vl_logic;
        o_riscv_de_immzeroextend_e: out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of width : constant is 1;
end riscv_de_ppreg;
