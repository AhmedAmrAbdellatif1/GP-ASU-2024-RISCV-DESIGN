package ranges;
    longint INT64_MAX = 64'h7FFFFFFFFFFFFFFF;
    longint INT64_MIN = 64'h8000000000000000;
    int     NO_TESTS  = 1000;
    int i;
    event failed;
    int counter=0;
endpackage